package types is

  subtype BYTE is std_logic_vector(7 downto 0);
  
end package types;
