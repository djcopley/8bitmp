package types is

  subtype REG_T is WORD;
  
end package types;
