package helpers is

  function my_func (L, R : std_logic) return std_logic;

end package;
