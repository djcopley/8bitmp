library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library cpu_lib;
use cpu_lib.helpers.all;

entity cpu is
  port(
    clk : in std_logic;
    rst : in std_logic
  );
end entity cpu;

architecture rtl of cpu is

begin

end architecture rtl;

