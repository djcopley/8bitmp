library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package constants is
  
  constant DATA_WIDTH : natural := 8;

end package constants;
